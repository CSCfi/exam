email.inspection.ready.subject=Tenttivastauksesi on arvioitu
email.inspection.new.subject=Sinut on lisätty arvioijaksi
email.enrolment.unit.pieces=kpl
email.enrolment.no.reservation=HUOM! tenttiakvaariota ei varattu
email.enrolment.no.enrolments=Ei ilmoittautuneita
email.weekly.report.subject=EXAM viikkokooste
email.machine.reservation.subject=Tenttitilavaraus
email.review.request.subject=Exam-tentti on annettu arvioitavaksesi
email.reservation.cancellation.subject=Tekemäsi varaus EXAM-tenttiin on peruttu
email.reservation.cancellation.info=Lisätietoja
email.template.inspection.done={0} on tehnyt oman osansa arvioinnista. Arviointi koskee tenttiä
email.template.inspection.comment=Arvioinnin palaute
email.template.link.to.review=Arviointiin
email.template.review.ready=Vastauksesi tenttiin {0} on arvioitu. Voit lukea alustavan arvioinnin ja palautteen täältä
email.template.main.system.info=Lopullisen arvosanan näet opintohallinnon järjestelmästä
email.template.inspector.new={0} on merkinnyt sinut arvioijaksi seuraavalle tentille
email.template.participation=Tentillä on {0} arvioitavaa suoritusta.
email.template.inspector.message=Saateviesti
email.template.link.to.exam=Tenttinäkymään
email.template.reservation.new=Olet varannut tenttipaikan tenttiakvaariosta. Tässä varauksesi tiedot
email.template.reservation.exam=Tentti: {0}
email.template.reservation.teacher=Opettaja: {0}
email.template.reservation.date=Tenttiaika: {0}
email.template.reservation.exam.duration=Tentin kesto: {0}
email.template.reservation.building=Rakennus: {0}
email.template.reservation.room=Luokka: {0}
email.template.reservation.machine=Kone: {0}
email.template.reservation.cancel.info=Peruthan ilmoittautumisesi, jos tenttisuunnitelmasi muuttuvat.
email.template.reservation.cancel.link.text=Varauksen peruminen
email.template.hello=Hei!
email.template.regards=Ystävällisin terveisin
email.template.admin=EXAM-ylläpito
email.template.reservation.cancel.message=Varauksesi EXAM-tenttiin {0} klo {1} tilassa {2} on jouduttu perumaan.
email.template.enrolment.first={0} kpl, joista ensimmäinen on tulossa {1}
email.template.weekly.report.enrolments=Ilmoittautumiset
email.template.weekly.report.enrolments.info=Opiskelijoita on ilmoittautunut tentteihisi seuraavasti
email.template.weekly.report.inspections=Arvioinnit
email.template.weekly.report.inspections.info=Sinulla on arvioimattomia vastauksia {0} kpl näissä tenteissä
