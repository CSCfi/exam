email.inspection.ready.subject=Ditt tentamenssvar är bedömt
email.inspection.comment.subject=Ny kommentar till bedömningen är tillsatt
email.enrolment.no.reservation=OBS! Du har inte ännu bokat tid för tentamen!
email.enrolment.no.enrolments=Inga bokningar
email.weekly.report.subject=Veckosammanfattning
email.machine.reservation.subject=Bokning av tentamenstid
email.machine.reservation.reminder.subject=Påminnelse om tentamensbokning
email.review.request.subject=Du är markerad som examinator för tentamen
email.reservation.cancellation.subject=Du har avbokat din tentamenstid
email.reservation.cancellation.subject.forced=Din bokning för tentamen "{0}" har avbokats
email.reservation.cancellation.info=Tilläggsinformation
email.template.inspection.done={0} har bedömt tentamen
email.template.inspection.comment=Meddelande till andra bedömare
email.template.link.to.review=Länk till återkoppling
email.template.review.ready=Din tentamen {0} är bedömd. Läs bedömningen här
email.template.review.autoevaluated=Bedömningen är automatisk och inte slutlig. Läraren kan vid behov ännu ändra bedömningen.
email.template.main.system.info=Kursens slutvitsord hittar du i studieregistret
email.template.inspector.new={0} har markerat dig som bedömare för tentamen
email.template.participation=Tentamen har {0} obedömda prestationer
email.template.inspector.message=Meddelandet
email.template.link.to.exam=Länk till tentamen
email.template.reservation.new=Du har bokat en tentamenstid. Här får du bokningsinformationen
email.template.reservation.exam=Tentamen: {0}
email.template.reservation.teacher=Ansvarslärare/Huvudansvarig tentator: {0}
email.template.reservation.date=Tid: {0}
email.template.reservation.exam.duration=Tentamens längd: {0}
email.template.reservation.building=Byggnad: {0}
email.template.reservation.room=Utrymme: {0}
email.template.reservation.machine=Dator: {0}
email.template.reservation.cancel.info=Kom ihåg att annullera din bokning om dina planer ändras!
email.template.reservation.cancel.link.text=Annullera bokningen
email.template.regards=Med vänliga hälsningar
email.template.admin=EXAM-administratörerna
email.template.reservation.cancel.message=Din bokning för tentamen {0} kl. {1} i {2} har avbokats
email.template.enrolment.first={0} st varav den första på {1}
email.template.weekly.report.enrolments=Bokningar
email.template.weekly.report.enrolments.info=Studerandena har bokat följande tider för dina tentamina
email.template.weekly.report.inspections=Obedömda prestationer
email.template.weekly.report.inspections.info=Du har {0} obedömda svar i följande tentamina
email.template.weekly.report.none=Det finns inga
email.template.reservation.cancel.message.student=Du har avbokat din tid till följande tentamen:
email.template.reservation.cancel.message.student.new.time=Du kan boka en ny tid till tentamen här
email.template.participant.notification.subject=Personlig tentamen {0}
email.template.participant.notification.title=En personlig tentamen är skapad för dig. Du bör boka tentamenstid i systemet.
email.template.participant.notification.title.examination.event=En personlig tentamen är skapad för dig. Du bör boka tentamenstid i EXAM systemet.
email.template.participant.notification.exam=Tentamen: {0}
email.template.participant.notification.teacher=Ansvarslärare/Tentator: {0}
email.template.participant.notification.exam.period=Tentamens giltighetstid: {0}
email.template.participant.notification.exam.event=Tillställning: {0}
email.template.participant.notification.exam.duration=Tentamens längd: {0} minuter
email.template.participant.notification.please.reserve=Boka tid.
email.template.reservation.new.student=Studerande {0} har bokat tid till personlig tentamen
email.template.exam.aborted.subject=Studerande har avbrutit sin personliga tentamen
email.template.exam.aborted.message=Studerande {0} har avbrutit sin personliga tentamen {1} och prestationen ska inte bedömas.
email.template.exam.returned.subject=En personlig tentamen är inlämnad
email.template.exam.returned.message=Studerande {0} har lämnat in sin personliga tentamen {1} för bedömning.
email.template.noshow.subject=Studerande kom inte till sin personliga tentamen, no-show
email.template.noshow.message=Studerande {0} har inte använt den tentamenstid som hen hade bokat för tentamen {1}, no-show.
ical.reservation.summary=Bokningen
ical.reservation.filename=bokning {0}
ical.reservation.room.info=Utrymme: {0}
email.template.language.inspection.subject=Språkgranskningen slutförd
email.template.language.inspection.approved=GODKÄND
email.template.language.inspection.rejected=UNDERKÄND
email.template.language.inspection.student=Studerande: {0}
email.template.language.inspection.done=Prestationen har genomgått språkgranskning med följande resultat.
email.template.language.inspection.statement.title=Utlåtande
email.template.language.inspection.result=Resultat: {0}
email.template.exam.returned.link=Länk till bedömningen
email.weekly.report.review.summary={0} tentamina (bedömning deadline {1})
email.template.maturity.participant.notification.subject=Ett mognadsprov har skapats för dig {0}
email.template.maturity.participant.notification.title=Ett mognadsprov har skapats för dig. Du måste boka tentamenstid i Exam.
email.template.maturity.exam.aborted.subject=Studerande har avbrutit mongadsprovet
email.template.maturity.exam.aborted.message=Studerande {0} har valt att avbryta mognadsprovet {1} och du skall inte bedöma prestationen.
email.template.maturity.exam.returned.subject=Mognadsprovet har inlämnats
email.template.maturity.exam.returned.message=Studerande {0} har utfört mognadsprov {1}
email.template.maturity.noshow.subject=Studerande kom inte till mognadsprovet (no show)
email.template.noshow.student.subject=Du kom inte till din bokade e-tentamen i EXAM
email.template.noshow.student.message=Du kom inte till din tentamen {0}{1} på din bokade tid.
email.template.reservation.change.subject=Tentamensdatorn utbytt: "{0}"
email.template.reservation.change.message=Hej, Exam-administratorn har bytt din tentamensdator till en annan dator.
email.template.reservation.change.previous=Föregående dator
email.template.reservation.change.current=Ny dator
email.template.reservation.exam.info=Information om tentamen
email.template.section.title=De sektioner du valt.
email.template.section.name=Namn
email.template.section.description=Beskrivning
email.examinationEvent.reminder.subject=Påminnelse om kommande tentamenstillfälle
email.examinationEvent.subject=Anmälan till tentamenstillfälle
email.examinationEvent.title=Du har anmält dig till ett tentamenstillfälle. Här är information om tentamenstillfället.
email.examinationEvent.date=Tentamenstillfället börjar: {0}
email.examinationEvent.file.info=I bilagan är en fil, men hjälp av vilket tentamen startas då tentamenstillfället har börjat.
email.examinationEvent.cancel.info=Du kommer ju ihåg att annullera din anmälan i tid, om dina planer ändrar!
email.examinationEvent.cancel.link.text=Ändring eller annullering av anmälan
email.examinationEvent.cancel.subject=Annullering av din anmälan
email.examinationEvent.cancel.message.student=Du har annullerat din anmälan till följande tentamenstillfälle:
email.examinationEvent.cancel.message.admin=Din anmälan till följande tentamenstillfälle har annullerats:
email.examinationEvent.cancel.message.student.new.time=Du kan anmäla dig på nytt till tentamenstillfället här.
clozeTest.blank.answer=blank
reports.scores.sectionScore=Poäng för ämnesområdet {0}
reports.scores.totalScore=Totala poäng i tentamen
reports.scores=Poäng
reports.studentFirstName=Förnamn
reports.studentLastName=Efternamn
reports.studentEmail=E-post
reports.studentId=Studentnummer
reports.question.type.essay=Essä
reports.question.type.cloze=Text med luckor
reports.question.type.multiplechoice=Flervalsfråga
reports.question.type.weightedmultiplechoide=Flervalsfråga
reports.question.type.claim=Påstående
reports.question=Fråga
