email.inspection.ready.subject=Ditt tentamenssvar är bedömt
email.inspection.comment.subject=Ny kommentar till bedömningen är tillsatt
email.enrolment.no.reservation=OBS! Du har inte ännu bokat tid för tentamen!
email.enrolment.no.enrolments=Inga bokningar
email.weekly.report.subject=Veckosammanfattning
email.machine.reservation.subject=Bokning
email.machine.reservation.reminder.subject = Påminnelse om bokning
email.review.request.subject=Du är markerad som examinator för tentamen
email.reservation.cancellation.subject=Bokningen du annulerar
email.reservation.cancellation.subject.forced=Din bokning för tentamen "{0}" är annulerad
email.reservation.cancellation.info=Tilläggsinformation
email.template.inspection.done={0} har bedömt tentamen
email.template.inspection.comment=Meddelande till andra bedömare
email.template.link.to.review=Länk till feedback
email.template.review.ready=Din tentamen {0} är bedömd. Läs den preliminära bedömningen här
email.template.review.autoevaluated=Bedömningen är automatisk och inte slutlig. Examinatorn kan vid behov ännu ändra den bedömningen.
email.template.main.system.info=Det slutliga vitsordet hittar du i studentregistret
email.template.inspector.new={0} har markerat dig som bedömare för tentamen
email.template.participation=Tentamen har {0} obedömda prestationer
email.template.inspector.message=Meddelandet
email.template.link.to.exam=Länk till tentamen
email.template.reservation.new=Du har bokat en tid. Här får du bokningens detaljer
email.template.reservation.exam=Tentamen: {0}
email.template.reservation.teacher=Ansvarslärare/Huvudansvarig tentator: {0}
email.template.reservation.date=Tid: {0}
email.template.reservation.exam.duration=Tentamens längd: {0}
email.template.reservation.building=Byggnad: {0}
email.template.reservation.room=Utrymme: {0}
email.template.reservation.machine=Dator: {0}
email.template.reservation.cancel.info=Kom ihåg att inhibera din bokning om dina planer ändras!
email.template.reservation.cancel.link.text=Inhibera bokningen
email.template.regards=Med vänliga hälsningar
email.template.admin=Systemadministratörerna
email.template.reservation.cancel.message=Din bokning för tentamen {0} kl. {1} i {2} har inhiberats
email.template.enrolment.first={0} st varav den första på {1}
email.template.weekly.report.enrolments=Bokningar
email.template.weekly.report.enrolments.info=Studerandena har bokat följande tider för dina tentamina
email.template.weekly.report.inspections=Obedömda prestationer
email.template.weekly.report.inspections.info=Du har {0} obedömda svar i följande tentamina
email.template.reservation.cancel.message.student=Du har inhiberat din tid till följande tentamen:
email.template.reservation.cancel.message.student.new.time=Du kan boka en ny tid till tentamen här
email.template.participant.notification.subject=Personlig tentamen {0}
email.template.participant.notification.title=En personlig tentamen är skapad för dig. Du bör boka tentamenstid i systemet.
email.template.participant.notification.exam=Tentamen: {0}
email.template.participant.notification.teacher=Ansvarslärare/Tentator: {0}
email.template.participant.notification.exam.period=Tentamens giltighetstid: {0}
email.template.participant.notification.exam.duration=Tentamens längd: {0} minuter
email.template.participant.notification.please.reserve=Boka tid.
email.template.reservation.new.student=Studerande {0} har bokat tid till personlig tentamen
email.template.exam.aborted.subject=Den personliga tentamen avbröts
email.template.exam.aborted.message=Studerande {0} har avbrutit tentamen {1}.
email.template.exam.returned.subject=Personliga tentamen är inlämnad
email.template.exam.returned.message=Studerande {0} har lämnat in sin personliga tentamen {1} för bedömning.
email.template.noshow.subject=Studerande {0} kom inte till sin personliga tentamen
email.template.noshow.message=Studerande {0} har inte använt bokad tid till tentamen {1}, no-show.
ical.reservation.summary=Bokningen
ical.reservation.filename=bokning {0}
ical.reservation.room.info=Utrymme: {0}
email.template.language.inspection.subject=Språkgranskningen slutförd
email.template.language.inspection.approved=GODKÄND
email.template.language.inspection.rejected=UNDERKÄND
email.template.language.inspection.student=Studerande: {0}
email.template.language.inspection.done=Prestationen har genomgått språkgranskning med följande resultat.
email.template.language.inspection.statement.title=Utlåtande
email.template.language.inspection.result=Resultat: {0}
email.template.exam.returned.link=Länk till bedömningen
email.weekly.report.review.summary={0} tentamina (bedömning deadline {1})
email.template.maturity.participant.notification.subject=Ett mognadsprov har skapats för dig {0}
email.template.maturity.participant.notification.title=Ett mognadsprov har skapats för dig. Du måste boka tentamenstid i Exam.
email.template.maturity.exam.aborted.subject=Studerande har avbrutit mongadsprovet
email.template.maturity.exam.aborted.message=Studerande {0} har valt att avbryta mognadsprovet {1} och du skall inte bedöma prestationen.
email.template.maturity.exam.returned.subject=Mognadsprovet har inlämnats
email.template.maturity.exam.returned.message=Studerande {0} har utfört mognadsprov {1}
email.template.maturity.noshow.subject=Studerande kom inte till mognadsprovet (no show)
email.template.noshow.student.subject=Et saapunut varaamaasi EXAM-tenttiin SV
email.template.noshow.student.message=Et saapunut tenttiin {0} ({1}) tenttivarauksen aikana. SV
