email.inspection.ready.subject=Ditt tentsvar är utvärderat
email.inspection.comment.subject=Ny kommentar på utvärdering
email.enrolment.no.reservation=OBS! Du har inte ännu bokat tid för tenten!
email.enrolment.no.enrolments=Inga tentbokningar
email.weekly.report.subject=Veckosammanfattning för dina tenter
email.machine.reservation.subject=Tentbokning
email.review.request.subject=Du har fått ett tentsvar för utvärdering
email.reservation.cancellation.subject=Din tentbokning är inhiberad
email.reservation.cancellation.info=Tilläggsinformation
email.template.inspection.done={0} har utvärderat sin del av tentsvaret som gäller tenten
email.template.inspection.comment=Feedback
email.template.link.to.review=Länk till feedback
email.template.review.ready=Ditt svar till tenten {0} är utvärderat. Läs den preliminära utvärderingen här
email.template.main.system.info=Det slutliga vitsordet hittar du i studentregistret
email.template.inspector.new={0} har markerat dig som utvärderare för tenten
email.template.participation=Tenten har {0} outvärderade svar
email.template.inspector.message=Meddelandet
email.template.link.to.exam=Länk till tenten
email.template.reservation.new=Du har bokat en tenttid. Här får du bokningens detaljer
email.template.reservation.exam=Tent: {0}
email.template.reservation.teacher=Tentator: {0}
email.template.reservation.date=Tenttid: {0}
email.template.reservation.exam.duration=Tentens längd: {0}
email.template.reservation.building=Byggnad: {0}
email.template.reservation.room=Klassrum: {0}
email.template.reservation.machine=Dator: {0}
email.template.reservation.cancel.info=Kom ihåg att inhibera din tentbokning om dina planer ändras!
email.template.reservation.cancel.link.text=Inhibera bokningen
email.template.regards=Mvh
email.template.admin=Systemadministratörerna
email.template.reservation.cancel.message=Din bokning för tenten {0} kl {1} i {2} har inhiberats
email.template.enrolment.first={0} st varav den första på {1}
email.template.weekly.report.enrolments=Tentbokningar
email.template.weekly.report.enrolments.info=Studerandena har bokat tider för dina tenter på följande sätt
email.template.weekly.report.inspections=Utvärderingar
email.template.weekly.report.inspections.info=Du har {0} outvärderade svar i följande tenter
email.template.reservation.cancel.message.student=Du har inhiberat din tid till följande tent:
email.template.reservation.cancel.message.student.new.time=Du kan boka en ny tid till tent
email.template.participant.notification.subject=Henkilökohtainen tentti {0} SV
email.template.participant.notification.title=Henkilökohtainen tentti on luotu. Opiskelijan tulee varata tenttiaika järjestelmästä. SV
email.template.participant.notification.exam=Tentti: {0} SV
email.template.participant.notification.teacher=Opettajat: {0} SV
email.template.participant.notification.exam.period=Tentin voimassaoloaika: {0} SV
email.template.participant.notification.exam.duration=Tentin kesto: {0} minuuttia SV
email.template.participant.notification.please.reserve=Varaa tenttiaika. SV
email.template.reservation.new.student=Opiskelija {0} on varannut tenttiajan henkilökohtaiseen tenttiin SV
email.template.exam.aborted.subject=Henkilökohtainen tentti on keskeytetty SV
email.template.exam.aborted.message=Opiskelija {0} on keskeyttänyt tentin {1}. SV
email.template.exam.returned.subject=Henkilökohtainen tentti on palautettu SV
email.template.exam.returned.message=Opiskelija {0} on palauttanut tentin {1} arvioitavaksi. SV
email.template.noshow.subject=Opiskelija ei saapunut henkilökohtaiseen tenttiin SV
email.template.noshow.message=Opiskelija {0} ei käyttänyt tenttiin {1} varaamaansa aikaa, no-show. SV

