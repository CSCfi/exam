email.inspection.ready.subject=Ditt tentsvar är utvärderat
email.inspection.new.subject=Du har fått tentator-rättigheter
email.enrolment.no.reservation=OBS! Du har inte ännu bokat tid i tentakvariet
email.enrolment.no.enrolments=Inga tentbokningar
email.weekly.report.subject=Exam-veckosammanfattning
email.machine.reservation.subject=Tentbokning
email.review.request.subject=Du har fått ett Exam-tentsvar för utvärdering
email.reservation.cancellation.subject=Din tentbokning är inhiberad
email.reservation.cancellation.info=Tilläggsinformation
email.template.inspection.done={0} har utvärderat sin del av tentsvaret som gäller tenten
email.template.inspection.comment=Feedback
email.template.link.to.review=Länk till feedback
email.template.review.ready=Ditt svar till tenten {0} är utvärderat. Läs den preliminära utvärderingen här
email.template.main.system.info=Det slutliga vitsordet hittar du i studentregistret
email.template.inspector.new={0} har markerat dig som utvärderare för tenten
email.template.participation=Tenten har {0} outvärderade svar
email.template.inspector.message=Meddelandet
email.template.link.to.exam=Länk till tenten
email.template.reservation.new=Du har bokat en tid i tentakvariet. Här får du bokningens detaljer
email.template.reservation.exam=Tent: {0}
email.template.reservation.teacher=Tentator: {0}
email.template.reservation.date=Tenttid: {0}
email.template.reservation.exam.duration=Tentens längd: {0}
email.template.reservation.building=Byggnad: {0}
email.template.reservation.room=Klassrum: {0}
email.template.reservation.machine=Dator: {0}
email.template.reservation.cancel.info=Kom ihåg att inhibera din tentbokning om dina planer ändras!
email.template.reservation.cancel.link.text=Inhibera bokningen
email.template.hello=Hej!
email.template.regards=Mvh
email.template.admin=EXAM-administratörerna
email.template.reservation.cancel.message=Din bokning för tenten {0} kl {1} i {2} har inhiberats
email.template.enrolment.first={0} st varav den första på {1}
email.template.weekly.report.enrolments=Tentboningar
email.template.weekly.report.enrolments.info=Studerandena har bokat tider för dina tenter på följande sätt
email.template.weekly.report.inspections=Utvärderingar
email.template.weekly.report.inspections.info=Du har {0} outvärderade svar kpl i följande tenter