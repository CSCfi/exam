email.inspection.ready.subject=Ditt tentsvar är utvärderat
email.inspection.comment.subject=Ny kommentar på utvärdering
email.enrolment.no.reservation=OBS! Du har inte ännu bokat tid för tenten!
email.enrolment.no.enrolments=Inga tentbokningar
email.weekly.report.subject=Veckosammanfattning för dina tenter
email.machine.reservation.subject=Tentbokning
email.review.request.subject=Du har fått ett tentsvar för utvärdering
email.reservation.cancellation.subject=Din tentbokning är inhiberad
email.reservation.cancellation.info=Tilläggsinformation
email.template.inspection.done={0} har utvärderat sin del av tentsvaret som gäller tenten
email.template.inspection.comment=Feedback
email.template.link.to.review=Länk till feedback
email.template.review.ready=Ditt svar till tenten {0} är utvärderat. Läs den preliminära utvärderingen här
email.template.main.system.info=Det slutliga vitsordet hittar du i studentregistret
email.template.inspector.new={0} har markerat dig som utvärderare för tenten
email.template.participation=Tenten har {0} outvärderade svar
email.template.inspector.message=Meddelandet
email.template.link.to.exam=Länk till tenten
email.template.reservation.new=Du har bokat en tenttid. Här får du bokningens detaljer
email.template.reservation.exam=Tent: {0}
email.template.reservation.teacher=Tentator: {0}
email.template.reservation.date=Tenttid: {0}
email.template.reservation.exam.duration=Tentens längd: {0}
email.template.reservation.building=Byggnad: {0}
email.template.reservation.room=Klassrum: {0}
email.template.reservation.machine=Dator: {0}
email.template.reservation.cancel.info=Kom ihåg att inhibera din tentbokning om dina planer ändras!
email.template.reservation.cancel.link.text=Inhibera bokningen
email.template.regards=Mvh
email.template.admin=Systemadministratörerna
email.template.reservation.cancel.message=Din bokning för tenten {0} kl {1} i {2} har inhiberats
email.template.enrolment.first={0} st varav den första på {1}
email.template.weekly.report.enrolments=Tentbokningar
email.template.weekly.report.enrolments.info=Studerandena har bokat tider för dina tenter på följande sätt
email.template.weekly.report.inspections=Utvärderingar
email.template.weekly.report.inspections.info=Du har {0} outvärderade svar i följande tenter
email.template.reservation.cancel.message.student=Du har inhiberat din tid till följande tent:
email.template.reservation.cancel.message.student.new.time=Du kan boka en ny tid till tent
email.template.participant.notification.subject=Personlig tent {0}
email.template.participant.notification.title=En personlig tent är skapad. Studeranden böra boka tenttid i systemet.
email.template.participant.notification.exam=Tent {0}
email.template.participant.notification.teacher=Lärare {0}
email.template.participant.notification.exam.period=Tentens giltighetstid {0}
email.template.participant.notification.exam.duration=Tenttid: {0} minuter
email.template.participant.notification.please.reserve=Boka tenttid.
email.template.reservation.new.student=Studerande {0} har bokat tid till personlig tent
email.template.exam.aborted.subject=Den personliga tenten avbröts
email.template.exam.aborted.message=Studerande {0} har avbrutit tenten {1}.
email.template.exam.returned.subject=Personliga tenten är inlämnad
email.template.exam.returned.message=Studerande {0} har lämnat in sin personlig tent {1} för utvärdering.
email.template.noshow.subject=Studerande {0} kom inte till sin personlig tent
email.template.noshow.message=Studerande {0} har inte använt bokad tid till tenten {1}, no-show.
ical.reservation.summary=Bokning
ical.reservation.filename=bokning{0}
ical.reservation.room.info=Tentutrymme: {0}
